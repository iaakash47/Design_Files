VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  LAYER LEF58_TYPE STRING ;
  LAYER LEF58_WIDTH STRING ;
END PROPERTYDEFINITIONS

UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.001 ;
LAYER NWELL
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
  PROPERTY LEF58_WIDTH "WIDTH 0.23 ;" ;
END NWELL

LAYER DIFF
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE DIFFUSION ;" ;
  PROPERTY LEF58_WIDTH "WIDTH 0.044 ;" ;
END DIFF

LAYER DIFF_18
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE DIFFUSION ;" ;
  PROPERTY LEF58_WIDTH "WIDTH 0.33 ;" ;
END DIFF_18

LAYER DIFF_25
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE DIFFUSION ;" ;
  PROPERTY LEF58_WIDTH "WIDTH 0.33 ;" ;
END DIFF_25

LAYER PIMP
  TYPE IMPLANT ;
  WIDTH 0.102 ;
  SPACING 0.17 ;
END PIMP

LAYER NIMP
  TYPE IMPLANT ;
  WIDTH 0.102 ;
  SPACING 0.17 ;
END NIMP

LAYER M1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.13 0.13 ;
  WIDTH 0.05 ;
  OFFSET 0.1 0.1 ;
  AREA 0.01 ;
  SPACING 0.05 ;
  WIREEXTENSION 0.105 ;
  MAXWIDTH 5 ;
  MINENCLOSEDAREA 0.2 ;
  RESISTANCE RPERSQ 0.1 ;
END M1

LAYER VIA1
  TYPE CUT ;
  SPACING 0.07 ;
  SPACING 0.07 LAYER M1 ;
  WIDTH 0.05 ;
  RESISTANCE 1.5 ;
END VIA1

LAYER M2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.164 0.164 ;
  WIDTH 0.056 ;
  OFFSET 0.15 0.15 ;
  AREA 0.016 ;
  SPACING 0.056 ;
  WIREEXTENSION 0.105 ;
  MAXWIDTH 5 ;
  MINENCLOSEDAREA 0.2 ;
  RESISTANCE RPERSQ 0.1 ;
END M2

LAYER VIA2
  TYPE CUT ;
  SPACING 0.07 ;
  SPACING 0.07 LAYER M2 ;
  WIDTH 0.05 ;
  RESISTANCE 1.5 ;
END VIA2

LAYER M3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.164 0.164 ;
  WIDTH 0.056 ;
  OFFSET 0.15 0.15 ;
  AREA 0.016 ;
  SPACING 0.056 ;
  WIREEXTENSION 0.105 ;
  MAXWIDTH 5 ;
  MINENCLOSEDAREA 0.2 ;
  RESISTANCE RPERSQ 0.1 ;
END M3

LAYER VIA3
  TYPE CUT ;
  SPACING 0.07 ;
  SPACING 0.07 LAYER M3 ;
  WIDTH 0.05 ;
  RESISTANCE 1.5 ;
END VIA3

LAYER M4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.164 0.164 ;
  WIDTH 0.056 ;
  OFFSET 0.15 0.15 ;
  AREA 0.016 ;
  SPACING 0.056 ;
  WIREEXTENSION 0.105 ;
  MAXWIDTH 5 ;
  MINENCLOSEDAREA 0.2 ;
  RESISTANCE RPERSQ 0.1 ;
END M4

LAYER VIA4
  TYPE CUT ;
  SPACING 0.07 ;
  SPACING 0.07 LAYER M4 ;
  WIDTH 0.05 ;
  RESISTANCE 1.5 ;
END VIA4

LAYER M5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.164 0.164 ;
  WIDTH 0.056 ;
  OFFSET 0.15 0.15 ;
  AREA 0.016 ;
  SPACING 0.056 ;
  MAXWIDTH 5 ;
  MINENCLOSEDAREA 0.2 ;
  RESISTANCE RPERSQ 0.1 ;
END M5

LAYER VIA5
  TYPE CUT ;
  SPACING 0.07 ;
  SPACING 0.07 LAYER M5 ;
  WIDTH 0.05 ;
  RESISTANCE 1.5 ;
END VIA5

LAYER M6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.164 0.164 ;
  WIDTH 0.056 ;
  OFFSET 0.15 0.15 ;
  AREA 0.016 ;
  SPACING 0.056 ;
  MAXWIDTH 5 ;
  MINENCLOSEDAREA 0.2 ;
  RESISTANCE RPERSQ 0.1 ;
END M6

LAYER VIA6
  TYPE CUT ;
  SPACING 0.07 ;
  SPACING 0.07 LAYER M6 ;
  WIDTH 0.05 ;
  RESISTANCE 1.5 ;
END VIA6

LAYER M7
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.164 0.164 ;
  WIDTH 0.056 ;
  OFFSET 0.15 0.15 ;
  AREA 0.016 ;
  SPACING 0.056 ;
  MAXWIDTH 5 ;
  MINENCLOSEDAREA 0.2 ;
  RESISTANCE RPERSQ 0.1 ;
END M7

LAYER M8
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.164 0.164 ;
  WIDTH 0.056 ;
  OFFSET 0.15 0.15 ;
  AREA 0.016 ;
  SPACING 0.056 ;
  MAXWIDTH 5 ;
  MINENCLOSEDAREA 0.2 ;
  RESISTANCE RPERSQ 0.1 ;
END M8

LAYER M9
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 1.74 1.74 ;
  WIDTH 0.16 ;
  OFFSET 0.15 0.15 ;
  AREA 0.055 ;
  SPACING 0.16 ;
  MAXWIDTH 10 ;
  MINENCLOSEDAREA 0.2 ;
  RESISTANCE RPERSQ 0.28 ;
END M9

LAYER MRDL
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 4.5 4.5 ;
  WIDTH 2 ;
  OFFSET 0.15 0.15 ;
  SPACING 2 ;
  MAXWIDTH 30 ;
  RESISTANCE RPERSQ 0.35 ;
END MRDL

LAYER VIARDL
  TYPE CUT ;
  SPACING 2 ;
  WIDTH 2 ;
  RESISTANCE 0.05 ;
END VIARDL

LAYER VIA7
  TYPE CUT ;
  SPACING 0.07 ;
  SPACING 0.08 LAYER M7 ;
  WIDTH 0.05 ;
  RESISTANCE 1.5 ;
END VIA7

LAYER VIA8
  TYPE CUT ;
  SPACING 0.12 ;
  SPACING 0.08 LAYER M8 ;
  WIDTH 0.13 ;
  RESISTANCE 0.1 ;
END VIA8

LAYER CO
  TYPE CUT ;
  SPACING 0.05 ;
  WIDTH 0.042 ;
END CO

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIARULE DIFFCON GENERATE DEFAULT
  LAYER DIFF ;
    ENCLOSURE 0.02 0.01 ;
  LAYER M1 ;
    ENCLOSURE 0.035 0.004 ;
  LAYER CO ;
    RECT -0.021 -0.021 0.021 0.021 ;
    SPACING 0.092 BY 0.092 ;
END DIFFCON

VIARULE DIFFCONC GENERATE
  LAYER DIFF ;
    ENCLOSURE 0.01 0.02 ;
  LAYER M1 ;
    ENCLOSURE 0.035 0.004 ;
  LAYER CO ;
    RECT -0.021 -0.021 0.021 0.021 ;
    SPACING 0.092 BY 0.092 ;
END DIFFCONC

VIARULE VIA12 GENERATE DEFAULT
  LAYER M1 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M2 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 1.500000 ;
END VIA12

VIARULE VIA12C GENERATE DEFAULT
  LAYER M1 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER M2 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 1.500000 ;
END VIA12C

VIARULE VIA12BAR GENERATE DEFAULT
  LAYER M1 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M2 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA1 ;
    RECT -0.025 -0.05 0.025 0.05 ;
    SPACING 0.135 BY 0.185 ;
    RESISTANCE 1.000000 ;
END VIA12BAR

VIARULE VIA12BARC GENERATE DEFAULT
  LAYER M1 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER M2 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA1 ;
    RECT -0.025 -0.05 0.025 0.05 ;
    SPACING 0.135 BY 0.185 ;
    RESISTANCE 1.000000 ;
END VIA12BARC

VIARULE VIA12LG GENERATE DEFAULT
  LAYER M1 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M2 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.185 BY 0.185 ;
    RESISTANCE 0.500000 ;
END VIA12LG

VIARULE VIA12LGC GENERATE DEFAULT
  LAYER M1 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER M2 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.185 BY 0.185 ;
    RESISTANCE 0.500000 ;
END VIA12LGC

VIARULE VIA23 GENERATE DEFAULT
  LAYER M2 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M3 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 1.500000 ;
END VIA23

VIARULE VIA23C GENERATE DEFAULT
  LAYER M2 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER M3 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 1.500000 ;
END VIA23C

VIARULE VIA23BAR GENERATE DEFAULT
  LAYER M2 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M3 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA2 ;
    RECT -0.025 -0.05 0.025 0.05 ;
    SPACING 0.135 BY 0.185 ;
    RESISTANCE 1.000000 ;
END VIA23BAR

VIARULE VIA23BARC GENERATE DEFAULT
  LAYER M2 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER M3 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA2 ;
    RECT -0.025 -0.05 0.025 0.05 ;
    SPACING 0.135 BY 0.185 ;
    RESISTANCE 1.000000 ;
END VIA23BARC

VIARULE VIA23LG GENERATE DEFAULT
  LAYER M2 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M3 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.185 BY 0.185 ;
    RESISTANCE 0.500000 ;
END VIA23LG

VIARULE VIA23LGC GENERATE DEFAULT
  LAYER M2 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER M3 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.185 BY 0.185 ;
    RESISTANCE 0.500000 ;
END VIA23LGC

VIARULE VIA34 GENERATE DEFAULT
  LAYER M3 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M4 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 1.500000 ;
END VIA34

VIARULE VIA34C GENERATE DEFAULT
  LAYER M3 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER M4 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 1.500000 ;
END VIA34C

VIARULE VIA34BAR GENERATE DEFAULT
  LAYER M3 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M4 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA3 ;
    RECT -0.025 -0.05 0.025 0.05 ;
    SPACING 0.135 BY 0.185 ;
    RESISTANCE 1.000000 ;
END VIA34BAR

VIARULE VIA34BARC GENERATE DEFAULT
  LAYER M3 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER M4 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA3 ;
    RECT -0.025 -0.05 0.025 0.05 ;
    SPACING 0.135 BY 0.185 ;
    RESISTANCE 1.000000 ;
END VIA34BARC

VIARULE VIA34LG GENERATE DEFAULT
  LAYER M3 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M4 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.185 BY 0.185 ;
    RESISTANCE 0.500000 ;
END VIA34LG

VIARULE VIA34LGC GENERATE DEFAULT
  LAYER M3 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER M4 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.185 BY 0.185 ;
    RESISTANCE 0.500000 ;
END VIA34LGC

VIARULE VIA45 GENERATE DEFAULT
  LAYER M4 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M5 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA4 ;
    RECT -0.025 -0.025 0.025 0.025 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 1.500000 ;
END VIA45

VIARULE VIA45C GENERATE
  LAYER M4 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER M5 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA4 ;
    RECT -0.025 -0.025 0.025 0.025 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 1.500000 ;
END VIA45C

VIARULE VIA45BAR GENERATE DEFAULT
  LAYER M4 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M5 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA4 ;
    RECT -0.025 -0.05 0.025 0.05 ;
    SPACING 0.135 BY 0.185 ;
    RESISTANCE 1.000000 ;
END VIA45BAR

VIARULE VIA45BARC GENERATE
  LAYER M4 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER M5 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA4 ;
    RECT -0.025 -0.05 0.025 0.05 ;
    SPACING 0.135 BY 0.185 ;
    RESISTANCE 1.000000 ;
END VIA45BARC

VIARULE VIA45LG GENERATE DEFAULT
  LAYER M4 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M5 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.185 BY 0.185 ;
    RESISTANCE 0.500000 ;
END VIA45LG

VIARULE VIA45LGC GENERATE
  LAYER M4 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER M5 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.185 BY 0.185 ;
    RESISTANCE 0.500000 ;
END VIA45LGC

VIARULE VIA56 GENERATE DEFAULT
  LAYER M5 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M6 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA5 ;
    RECT -0.025 -0.025 0.025 0.025 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 1.500000 ;
END VIA56

VIARULE VIA56C GENERATE
  LAYER M5 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER M6 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA5 ;
    RECT -0.025 -0.025 0.025 0.025 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 1.500000 ;
END VIA56C

VIARULE VIA56BAR GENERATE DEFAULT
  LAYER M5 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M6 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA5 ;
    RECT -0.025 -0.05 0.025 0.05 ;
    SPACING 0.135 BY 0.185 ;
    RESISTANCE 1.000000 ;
END VIA56BAR

VIARULE VIA56BARC GENERATE
  LAYER M5 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER M6 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA5 ;
    RECT -0.025 -0.05 0.025 0.05 ;
    SPACING 0.135 BY 0.185 ;
    RESISTANCE 1.000000 ;
END VIA56BARC

VIARULE VIA56LG GENERATE DEFAULT
  LAYER M5 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M6 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.185 BY 0.185 ;
    RESISTANCE 0.500000 ;
END VIA56LG

VIARULE VIA56LGC GENERATE
  LAYER M5 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER M6 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.185 BY 0.185 ;
    RESISTANCE 0.500000 ;
END VIA56LGC

VIARULE VIA67 GENERATE DEFAULT
  LAYER M6 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M7 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA6 ;
    RECT -0.025 -0.025 0.025 0.025 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 1.500000 ;
END VIA67

VIARULE VIA67C GENERATE
  LAYER M6 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER M7 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA6 ;
    RECT -0.025 -0.025 0.025 0.025 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 1.500000 ;
END VIA67C

VIARULE VIA67BAR GENERATE DEFAULT
  LAYER M6 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M7 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA6 ;
    RECT -0.025 -0.05 0.025 0.05 ;
    SPACING 0.135 BY 0.185 ;
    RESISTANCE 1.000000 ;
END VIA67BAR

VIARULE VIA67BARC GENERATE
  LAYER M6 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER M7 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA6 ;
    RECT -0.025 -0.05 0.025 0.05 ;
    SPACING 0.135 BY 0.185 ;
    RESISTANCE 1.000000 ;
END VIA67BARC

VIARULE VIA67LG GENERATE DEFAULT
  LAYER M6 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M7 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA6 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.185 BY 0.185 ;
    RESISTANCE 0.500000 ;
END VIA67LG

VIARULE VIA67LGC GENERATE
  LAYER M6 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER M7 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA6 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.185 BY 0.185 ;
    RESISTANCE 0.500000 ;
END VIA67LGC

VIARULE VIA78 GENERATE DEFAULT
  LAYER M7 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M8 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA7 ;
    RECT -0.025 -0.025 0.025 0.025 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 1.500000 ;
END VIA78

VIARULE VIA78C GENERATE
  LAYER M7 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER M8 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA7 ;
    RECT -0.025 -0.025 0.025 0.025 ;
    SPACING 0.12 BY 0.12 ;
    RESISTANCE 1.500000 ;
END VIA78C

VIARULE VIA78BAR GENERATE DEFAULT
  LAYER M7 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M8 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA7 ;
    RECT -0.025 -0.05 0.025 0.05 ;
    SPACING 0.135 BY 0.185 ;
    RESISTANCE 1.000000 ;
END VIA78BAR

VIARULE VIA78BARC GENERATE
  LAYER M7 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER M8 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA7 ;
    RECT -0.025 -0.05 0.025 0.05 ;
    SPACING 0.135 BY 0.185 ;
    RESISTANCE 1.000000 ;
END VIA78BARC

VIARULE VIA78LG GENERATE DEFAULT
  LAYER M7 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER M8 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA7 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.185 BY 0.185 ;
    RESISTANCE 0.500000 ;
END VIA78LG

VIARULE VIA78LGC GENERATE
  LAYER M7 ;
    ENCLOSURE 0.005 0.03 ;
  LAYER M8 ;
    ENCLOSURE 0.03 0.005 ;
  LAYER VIA7 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.185 BY 0.185 ;
    RESISTANCE 0.500000 ;
END VIA78LGC

VIARULE VIA89 GENERATE DEFAULT
  LAYER M8 ;
    ENCLOSURE 0.03 0.015 ;
  LAYER M9 ;
    ENCLOSURE 0.03 0.015 ;
  LAYER VIA8 ;
    RECT -0.065 -0.065 0.065 0.065 ;
    SPACING 0.25 BY 0.25 ;
    RESISTANCE 0.100000 ;
END VIA89

VIARULE VIA89C GENERATE
  LAYER M8 ;
    ENCLOSURE 0.015 0.03 ;
  LAYER M9 ;
    ENCLOSURE 0.03 0.015 ;
  LAYER VIA8 ;
    RECT -0.065 -0.065 0.065 0.065 ;
    SPACING 0.25 BY 0.25 ;
    RESISTANCE 0.100000 ;
END VIA89C

VIARULE VIARDL GENERATE
  LAYER M9 ;
    ENCLOSURE 0.05 0.05 ;
  LAYER MRDL ;
    ENCLOSURE 0.05 0.05 ;
  LAYER VIARDL ;
    RECT -1 -1 1 1 ;
    SPACING 4 BY 4 ;
    RESISTANCE 0.050000 ;
END VIARDL

MACRO PLL
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 113.223 BY 48.108 ;
  SYMMETRY X Y R90 ;
 

  PIN Vss
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 16.062 -6.38 16.112 -6.33 ;
    END
  END Vss
  PIN Vout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.13 -3.264 21.18 -3.214 ;
    END
  END Vout
  PIN Vdd
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 6.22 0.266 6.276 0.322 ;
    END
  END Vdd
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M2 ;
        RECT 2.724 -7.53 2.78 -7.474 ;
    END
  END gnd!
  PIN Vref
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0 -1.08 0.05 -1.03 ;
    END
  END Vref
  OBS
    LAYER DIFF ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER DIFF_18 ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER PO ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER M1 ;
      POLYGON -2.963 -16.427 -2.963 1.547 23.139 1.547 23.139 -0.98 -0.05 -0.98 -0.05 -1.13 0.1 -1.13 0.1 -0.98 23.139 -0.98 23.139 -6.28 16.012 -6.28 16.012 -6.43 16.162 -6.43 16.162 -6.28 23.139 -6.28 23.139 -16.427 ;
    LAYER VIA1 ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER M2 ;
      POLYGON -2.963 -16.427 -2.963 1.547 23.139 1.547 23.139 0.378 6.164 0.378 6.164 0.21 6.332 0.21 6.332 0.378 23.139 0.378 23.139 -3.158 21.074 -3.158 21.074 -3.32 21.236 -3.32 21.236 -3.158 23.139 -3.158 23.139 -7.418 2.668 -7.418 2.668 -7.586 2.836 -7.586 2.836 -7.418 23.139 -7.418 23.139 -16.427 ;
    LAYER VIA2 ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER M3 ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER VIA3 ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER M4 ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER VIA4 ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER M5 ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER VIA5 ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER M6 ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER VIA6 ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER M7 ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER VIA7 ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER M8 ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER VIA8 ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER M9 ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER CO ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER M1PIN ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER M2PIN ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER M3PIN ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER M4PIN ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER M5PIN ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER M6PIN ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER M7PIN ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER M8PIN ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER M9PIN ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER MRDL ;
      RECT -2.963 -16.427 23.139 1.547 ;
    LAYER VIARDL ;
      RECT -2.963 -16.427 23.139 1.547 ;
  END
END PLL

END LIBRARY
